-- Package Declaration Section
package pixel_bus is
   
end package pixel_bus;
 
-- Package Body Section
package body pixel_bus is
 
end package body pixel_bus;