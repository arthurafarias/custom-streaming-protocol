-- Package Declaration Section
package custom_stream is
   
end package custom_stream;
 
-- Package Body Section
package body custom_stream is
 
end package body custom_stream;