entity pixel_bus_split_1x2_tb is
end pixel_bus_split_1x2_tb;

architecture impl of pixel_bus_split_1x2_tb is
begin
end impl;