entity pixel_bus_concat
end pixel_bus_concat;

architecture impl of pixel_bus_concat is
begin
end impl;