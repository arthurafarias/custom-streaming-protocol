entity custom_stream_passthrough is
-- generic();
-- port();
end custom_stream_passthrough;

architecture impl of custom_stream_passthrough is
begin
    
end impl;