entity pixel_bus_passthrough is
-- generic();
-- port();
end pixel_bus_passthrough;

architecture impl of pixel_bus_passthrough is
begin
    
end impl;