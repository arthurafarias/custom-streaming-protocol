entity pixel_bus_inspect is
-- generic();
-- port();
end pixel_bus_inspect;

architecture impl of pixel_bus_inspect is
begin
end impl;