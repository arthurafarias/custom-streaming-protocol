entity custom_stream_product_cross is
-- generic();
-- port();
end custom_stream_product_cross;

architecture impl of custom_stream_product_cross is
begin
    
end impl;